module ProgramCounter (
	input			clk,
	input			
);
