module InstrDec (
	input				clk,
	input [6:0] opcode,
	input	[6:0] 
);
